// jtag_to_pio_pd.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module jtag_to_pio_pd (
		input  wire       clk_i_clk,       //   clk_i.clk
		output wire [7:0] pio_o_export,    //   pio_o.export
		input  wire       reset_i_reset_n  // reset_i.reset_n
	);

	wire  [31:0] master_0_master_readdata;              // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;           // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;               // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                  // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;            // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;         // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                 // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;             // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire         mm_interconnect_0_pio_0_s1_chipselect; // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;   // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;    // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;      // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;  // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata

	jtag_to_pio_pd_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_i_clk),                     //          clk.clk
		.clk_reset_reset      (~reset_i_reset_n),              //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	jtag_to_pio_pd_pio_0 pio_0 (
		.clk        (clk_i_clk),                             //                 clk.clk
		.reset_n    (reset_i_reset_n),                       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (pio_o_export)                           // external_connection.export
	);

	jtag_to_pio_pd_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_i_clk),                             //                                clk_0_clk.clk
		.master_0_clk_reset_reset_bridge_in_reset_reset (~reset_i_reset_n),                      // master_0_clk_reset_reset_bridge_in_reset.reset
		.pio_0_reset_reset_bridge_in_reset_reset        (~reset_i_reset_n),                      //        pio_0_reset_reset_bridge_in_reset.reset
		.master_0_master_address                        (master_0_master_address),               //                          master_0_master.address
		.master_0_master_waitrequest                    (master_0_master_waitrequest),           //                                         .waitrequest
		.master_0_master_byteenable                     (master_0_master_byteenable),            //                                         .byteenable
		.master_0_master_read                           (master_0_master_read),                  //                                         .read
		.master_0_master_readdata                       (master_0_master_readdata),              //                                         .readdata
		.master_0_master_readdatavalid                  (master_0_master_readdatavalid),         //                                         .readdatavalid
		.master_0_master_write                          (master_0_master_write),                 //                                         .write
		.master_0_master_writedata                      (master_0_master_writedata),             //                                         .writedata
		.pio_0_s1_address                               (mm_interconnect_0_pio_0_s1_address),    //                                 pio_0_s1.address
		.pio_0_s1_write                                 (mm_interconnect_0_pio_0_s1_write),      //                                         .write
		.pio_0_s1_readdata                              (mm_interconnect_0_pio_0_s1_readdata),   //                                         .readdata
		.pio_0_s1_writedata                             (mm_interconnect_0_pio_0_s1_writedata),  //                                         .writedata
		.pio_0_s1_chipselect                            (mm_interconnect_0_pio_0_s1_chipselect)  //                                         .chipselect
	);

endmodule
