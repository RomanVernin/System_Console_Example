
module jtag_to_pio_pd (
	clk_i_clk,
	pio_o_export,
	reset_i_reset_n);	

	input		clk_i_clk;
	output	[7:0]	pio_o_export;
	input		reset_i_reset_n;
endmodule
